/*
	This file implements the instruction fetch stage of ARVI's datapath.
*/

`include "arvi_defines.svh"
