`ifndef __DEFINES
`define __DEFINES
//`define SIMULATION

`define INSTRUCTION_SIZE 31
`define WORD_SIZE 31
`define XLEN 32
// Start address
`define PC_RESET 32'h80000000

`define PROGRAM_DATA "./test/asm/addi.bin"

// Extensions
//`define __ATOMIC

`endif
