`timescale 1ns / 1ps

module BRIDGE_2X1(
	input i_clk,
	input i_rst


	);

endmodule