import "DPI-C" function void new_instruction (input int inst);