`ifndef __M_INSTRUCTIONS
`define __M_INSTRUCTIONS

`define MUL    3'b000
`define MULH   3'b001
`define MULHSU 3'b010
`define MULHU  3'b011
`define DIV    3'b100
`define DIVU   3'b101
`define REM    3'b110
`define REMU   3'b111

`endif