`ifndef __ATOMIC_INSTRUCTIONS
`define __ATOMIC_INSTRUCTIONS

`define LR 		5'b00010
`define SC 		5'b00011
`define AMOSWAP 5'b00001
`define AMOADD  5'b00000
`define AMOXOR  5'b00100
`define AMOAND  5'b01100
`define AMOOR   5'b01000
`define AMOMIN  5'b10000
`define AMOMAX  5'b10100
`define AMOMINU 5'b11000
`define AMOMAXU 5'b11100

`endif