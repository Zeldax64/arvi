import "DPI-C" function void new_instruction (input int inst, input int cycles);