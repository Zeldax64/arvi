`ifdef __ATOMIC



`endif